`timescale 1ns / 1ps

module buffer(
	input a,
	output y
);

assign y=a;

endmodule